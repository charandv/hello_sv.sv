module hello_sv;
  initial begin
    $display("Hello DV World!");
  end
endmodule
